**.subckt untitled vg vd
*.opin vg
*.opin vd
XM1 vd vg GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
v1 vg GND 0
v2 vd GND 0.9
**** begin user architecture code

.option TEMP=27C
.option dccap post brief accurate nomod

.dc v1 0 3 0.01

.control
  run
  plot (-i(v2))
.endc

.save all


 ** manual skywater pdks install (with patches applied)
* .lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param mc_mm_switch=0
.param mc_pr_switch=0

**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
