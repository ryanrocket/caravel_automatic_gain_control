**.subckt test_nmos G1v8 D1v8 B
*.ipin G1v8
*.ipin D1v8
*.ipin B
Vd1 D1v8 net1 0
Vd3 D3v3 net2 0
Vd2 D1v8 net3 0
Vd4 D5v0 net4 0
E1 D5v0 0 D1v8 0 '5/1.8' 
E2 D3v3 0 D1v8 0 '3.3/1.8' 
E3 G5v0 0 G1v8 0 '5/1.8' 
E4 G3v3 0 G1v8 0 '3.3/1.8' 
Vd5 D10v5 net5 0
E5 D10v5 0 D1v8 0 '10.5/1.8' 
E6 D16v0 0 D1v8 0 '16.0/1.8' 
Vd6 D16v0 net6 0
Vd7 D1v8 net7 0
E7 D20v0 0 D1v8 0 '20.0/1.8' 
XM1 net1 G1v8 S B sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 net3 G1v8 S B sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net2 G3v3 S B sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 net4 G5v0 S B sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 net5 G5v0 S B sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 net6 G5v0 S B sky130_fd_pr__nfet_g5v0d16v0 L=0.7 W=5.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
Vd8 D1v8 net8 0
XM7 net7 G1v8 S B sky130_fd_pr__nfet_20v0 L=2.95 W=29.41 m=1
XM16 net8 G1v8 S B sky130_fd_pr__nfet_20v0_zvt W=30 L=5 m=1
**** begin user architecture code

* this experimental option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1
.option savecurrents
vg G1v8 0 1.8
vs s 0 0
vd D1v8 0 1.8
vb b 0 0
.control
save all
dc vd 0 1.8 0.01 vg 0 1.8 0.2
* dc vd 0 1.8 0.01 vg 0 1.2 0.1
plot all.vd1#branch vs D1v8
*plot all.vd2#branch vs D1v8
plot all.vd3#branch vs D3v3
*plot all.vd4#branch vs D5v0
plot all.vd5#branch vs D10v5
*plot all.vd6#branch vs D16v0
plot all.vd8#branch vs D1v8
plot all.vd7#branch vs D1v8
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
op
write test_nmos.raw
.endc



** manual skywater-pdk install (with patches applied).

** opencircuitdesign pdks install

 ** manual skywater pdks install (with patches applied)
* .lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param mc_mm_switch=0
.param mc_pr_switch=0

**** end user architecture code
**.ends
** flattened .save nodes
.save I(Vd1)
.save I(Vd3)
.save I(Vd2)
.save I(Vd4)
.save I(Vd5)
.save I(Vd6)
.save I(Vd7)
.save I(Vd8)
.end
