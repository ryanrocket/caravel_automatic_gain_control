** sch_path:
*+ /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/user_analog_project_wrapper.sch
**.subckt user_analog_project_wrapper in1 in2 vdd1 gnd1 dsa_ctr1 dsa_ctr2 dsa_ctr3 dsa_ctr4 pd_out
*+ out1 out2 gnd2 gnd3 gnd4 vdd2 vdd3 vdd4
*.ipin in1
*.ipin in2
*.ipin vdd1
*.ipin gnd1
*.ipin dsa_ctr1
*.ipin dsa_ctr2
*.ipin dsa_ctr3
*.ipin dsa_ctr4
*.opin pd_out
*.opin out1
*.opin out2
*.ipin gnd2
*.ipin gnd3
*.ipin gnd4
*.ipin vdd2
*.ipin vdd3
*.ipin vdd4
XDSA1 dsa_ctr1 dsa_ctr2 dsa_ctr3 dsa_ctr4 in2 vdd3 gnd3 net2 dsa
XDSA2 dsa_ctr1 dsa_ctr2 dsa_ctr3 dsa_ctr4 in1 vdd4 gnd4 net1 dsa
XLNA1 vdd2 vdd2 net1 net2 out1 out2 gnd2 gnd2 cmfb-negfb-revision
X1 out1 out2 net3 vdd1 pd_out gnd1 balaced-pd
R7 vdd2 net3 sky130_fd_pr__res_generic_po W=1 L=1 m=1
R1 net3 gnd1 sky130_fd_pr__res_generic_po W=1 L=1 m=1
**** begin user architecture code
?
**** end user architecture code
**.ends

* expanding   symbol:  /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/dsa.sym
*+ # of pins=8
** sym_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/dsa.sym
** sch_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/dsa.sch
.subckt dsa  ctr1 ctr2 ctr3 ctr4 in vdd gnd out
*.ipin in
*.ipin gnd
*.ipin vdd
*.ipin ctr1
*.ipin ctr2
*.ipin ctr3
*.ipin ctr4
*.opin out
XSPDT1 in ctr1 net1 net2 gnd vdd spdt
XSPDT2 net2 ctr2 net3 net4 gnd vdd spdt
XSPDT3 net4 ctr3 net5 net6 gnd vdd spdt
XSPDT4 net6 ctr4 net7 out gnd vdd spdt
XR1 net1 net2 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1 mult=1 m=1
XR2 net4 net3 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1 mult=1 m=1
XR3 net5 net6 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1 mult=1 m=1
XR4 net7 out gnd sky130_fd_pr__res_xhigh_po_0p35 L=1 mult=1 m=1
.ends


* expanding   symbol:
*+  /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/lownoiseamplifier/cmfb-negfb-revision.sym # of pins=8
** sym_path:
*+ /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/lownoiseamplifier/cmfb-negfb-revision.sym
** sch_path:
*+ /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/lownoiseamplifier/cmfb-negfb-revision.sch
.subckt cmfb-negfb-revision  vdd1 vdd2 in1 in2 out1 out2 gnd1 gnd2
*.ipin gnd1
*.ipin gnd2
*.ipin vdd1
*.ipin vdd2
*.ipin in1
*.ipin in2
*.opin out1
*.opin out2
XM1 out1 in1 net1 gnd1 sky130_fd_pr__nfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out2 in2 net1 gnd1 sky130_fd_pr__nfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 net2 gnd2 gnd2 sky130_fd_pr__nfet_01v8 L=0.15 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 net2 gnd2 gnd2 sky130_fd_pr__nfet_01v8 L=0.15 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 out1 net3 vdd2 vdd2 sky130_fd_pr__pfet_01v8 L=0.15 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 out2 net3 vdd2 vdd2 sky130_fd_pr__pfet_01v8 L=0.15 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R7 vdd1 net2 sky130_fd_pr__res_generic_po W=1 L=1 m=1
XR8 out2 net3 gnd1 sky130_fd_pr__res_high_po_0p35 L=1 mult=1 m=1
XR1 net3 out1 gnd1 sky130_fd_pr__res_high_po_0p35 L=1 mult=1 m=1
.ends


* expanding   symbol:
*+  /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/powerdetector/balaced-pd.sym # of pins=6
** sym_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/powerdetector/balaced-pd.sym
** sch_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/powerdetector/balaced-pd.sch
.subckt balaced-pd  in1 in2 vbias vdd output gnd
*.ipin vdd
*.ipin gnd
*.opin output
*.ipin in1
*.ipin in2
*.ipin vbias
XM11 output net3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net3 net2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 net2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 vbias gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net1 in1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 net1 in2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 net3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net1 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/spdt.sym
*+ # of pins=6
** sym_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/spdt.sym
** sch_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/spdt.sch
.subckt spdt  in ctr out1 out2 gnd vdd
*.ipin in
*.ipin ctr
*.ipin gnd
*.ipin vdd
*.opin out1
*.opin out2
XINV1 vdd ctr gnd net1 inverter
XTG1 vdd ctr in gnd net1 out1 transgate
XTG2 vdd net1 in gnd ctr out2 transgate
XINV1 vdd ctr gnd net1 inverter
.ends


* expanding   symbol:
*+  /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/inverter.sym # of pins=4
** sym_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/inverter.sym
** sch_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/inverter.sch
.subckt inverter  vdd in gnd out
*.ipin in
*.ipin gnd
*.ipin vdd
*.opin out
XM1 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/transgate.sym # of pins=6
** sym_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/transgate.sym
** sch_path: /Volumes/WORK_DRIVE/caravel_automatic_gain_control/xschem/attenuator/transgate.sch
.subckt transgate  vdd ctr2 in gnd ctr1 out
*.ipin in
*.ipin ctr2
*.ipin ctr1
*.ipin vdd
*.ipin gnd
*.opin out
XM1 in ctr1 out gnd sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 in ctr2 out vdd sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
