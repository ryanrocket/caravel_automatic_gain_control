**.subckt dsa cntrl1 cntrl2 cntrl3 cntrl4 in out gnd vbias vdd
*.ipin cntrl1
*.ipin cntrl2
*.ipin cntrl3
*.ipin cntrl4
*.ipin in
*.opin out
*.ipin gnd
*.ipin vbias
*.ipin vdd
R1 net1 net2 50 m=1
R2 net3 net4 200 m=1
XDTG1 in cntrl1 vdd vbias gnd net2 net1 transgate-full
XDTG2 net2 cntrl2 vdd vbias gnd net4 net3 transgate-full
R3 net5 net6 1k m=1
XDTG3 net4 cntrl3 vdd vbias gnd net6 net5 transgate-full
R4 net7 out 10k m=1
XDTG4 net6 cntrl4 vdd vbias gnd out net7 transgate-full
**** begin user architecture code
 ** manual skywater pdks install (with patches applied)
* .lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param mc_mm_switch=0
.param mc_pr_switch=0



.tran 0.000001s 0.0001s
.save all


**** end user architecture code
**.ends

* expanding   symbol:  transgate-full.sym # of pins=7
* sym_path: /home/u5921_ryanwan/design/FB1/xschem/transgate-full.sym
* sch_path: /home/u5921_ryanwan/design/FB1/xschem/transgate-full.sch
.subckt transgate-full  in cntrl vdd vbias gnd out2 out1
*.ipin cntrl
*.ipin vdd
*.ipin in
*.ipin gnd
*.ipin vbias
*.opin out2
*.opin out1
XI1 vdd gnd net1 cntrl basic-invert
XTG1 in out1 gnd vbias net1 cntrl gate-switch
XTG2 in out2 gnd vbias cntrl net1 gate-switch
.ends


* expanding   symbol:  basic-invert.sym # of pins=4
* sym_path: /home/u5921_ryanwan/design/FB1/xschem/basic-invert.sym
* sch_path: /home/u5921_ryanwan/design/FB1/xschem/basic-invert.sch
.subckt basic-invert  vdd gnd out in
*.ipin in
*.ipin gnd
*.ipin vdd
*.opin out
XM1 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  gate-switch.sym # of pins=6
* sym_path: /home/u5921_ryanwan/design/FB1/xschem/gate-switch.sym
* sch_path: /home/u5921_ryanwan/design/FB1/xschem/gate-switch.sch
.subckt gate-switch  in out gnd vbias cntrl2 cntrl1
*.ipin in
*.ipin vbias
*.ipin gnd
*.opin out
*.ipin cntrl1
*.ipin cntrl2
XM5 in cntrl2 out vbias sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 out cntrl1 in gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

** flattened .save nodes
.end
