**.subckt n_diffamp PLUS MINUS OUT NBIAS
*.ipin PLUS
*.ipin MINUS
*.opin OUT
*.ipin NBIAS
XM1 net1 PLUS S GND sky130_fd_pr__nfet_01v8_lvt L=0.3 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 OUT MINUS S GND sky130_fd_pr__nfet_01v8_lvt L=0.3 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 OUT net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.8 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 net1 net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.8 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 net2 NBIAS GND GND sky130_fd_pr__nfet_01v8 L=1.2 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XR1 GND S GND sky130_fd_pr__res_xhigh_po_0p35 L=50 mult=1 m=1
V1 PLUS GND 0.7
V2 NBIAS GND 0.9
V3 VDD GND 1.8
V4 MINUS GND 0.7
V5 S net2 0
**** begin user architecture code

.lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* Mismatch parameters
* Resistor/ef/tech/SW.2/sky130A/libs.tech/ngspice/Capacitor
* Special cells
* All models
* Corner

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
**** begin user architecture code

.options savecurrents
.control
save @m.xm5.msky130_fd_pr__nfet_01v8[gm]
save all
op
write n_diffamp.raw
.endc


**** end user architecture code
** flattened .save nodes
.end
