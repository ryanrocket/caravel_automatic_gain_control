**.subckt cs-exper
XM1 drain gate source GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
V1 net1 GND SIN(0 0.3 40)
C1 gate net1 500u m=1
R1 gate GND 1k m=1
R2 net3 gate 880 m=1
R3 source GND 1k m=1
R4 net2 drain 45k m=1
V2 net2 GND 1.8
V3 net3 GND 1.8
C2 source GND 500u m=1
**** begin user architecture code
 ** manual skywater pdks install (with patches applied)
* .lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param mc_mm_switch=0
.param mc_pr_switch=0



.tran 0.001s 0.1s
.control
  run
  plot v(drain) v(gate) v(source)
  plot -i(v2)
.endc
.save all


**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
