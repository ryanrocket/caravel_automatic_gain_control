**.subckt test_res P M B
*.ipin P
*.ipin M
*.ipin B
XR1 M net1 B sky130_fd_pr__res_iso_pw W=2.65 L=2.65 mult=1 m=1
Vr1 P net1 0
Vr2 P net2 0
R2 M net2 B sky130_fd_pr__res_generic_nd W=1 L=1 mult=1 m=1
Vr3 P net3 0
R3 M net3 B sky130_fd_pr__res_generic_pd W=1 L=1 mult=1 m=1
Vr4 P net4 0
R4 M net4 sky130_fd_pr__res_generic_po W=1 L=1 mult=1 m=1
Vr5 P net5 0
XR5 M net5 B sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
Vr6 P net6 0
XR6 M net6 B sky130_fd_pr__res_high_po_0p35 L=1 mult=1 m=1
Vr7 P net7 0
XR7 M net7 B sky130_fd_pr__res_high_po_0p69 L=0.69 mult=1 m=1
Vr8 P net8 0
XR8 M net8 B sky130_fd_pr__res_high_po_1p41 L=1.41 mult=1 m=1
Vr9 P net9 0
XR9 M net9 B sky130_fd_pr__res_xhigh_po W=1 L=1 mult=1 m=1
Vr10 P net10 0
XR10 M net10 B sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
Vr11 P net11 0
XR11 M net11 B sky130_fd_pr__res_xhigh_po_0p69 L=0.69 mult=1 m=1
Vr12 P net12 0
XR12 M net12 B sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
**** begin user architecture code


vp P 0 1.8
vm M 0 0
vb B 0 0
.control
save all
* dc vp 0 3 0.01
dc temp -40 140 1
*plot v(p,m) / vr1#branch
*plot v(p,m) / vr2#branch
*plot v(p,m) / vr3#branch
plot v(p,m) / vr4#branch
plot v(p,m) / vr5#branch
plot v(p,m) / vr6#branch
*plot v(p,m) / vr7#branch
*plot v(p,m) / vr8#branch
plot v(p,m) / vr9#branch
plot v(p,m) / vr10#branch
*plot v(p,m) / vr11#branch
*plot v(p,m) / vr12#branch

.endc


 ** manual skywater pdks install (with patches applied)
* .lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param mc_mm_switch=0
.param mc_pr_switch=0

**** end user architecture code
**.ends
** flattened .save nodes
.save I(Vr1)
.save I(Vr2)
.save I(Vr3)
.save I(Vr4)
.save I(Vr5)
.save I(Vr6)
.save I(Vr7)
.save I(Vr8)
.save I(Vr9)
.save I(Vr10)
.save I(Vr11)
.save I(Vr12)
.end
