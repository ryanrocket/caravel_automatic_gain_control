**.subckt FB1 vg vd
*.opin vg
*.opin vd
XM1 vd vg GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
v1 vg GND 1
v2 vd GND 0
**** begin user architecture code

.option TEMP=27C

.dc v2 0 3 0.01

.control
  set color0 = rgb:f/f/f
  alter @v1[dc] = 1
  print @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
  run
  alter @v1[dc] = 1.2
  print @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
  run
  alter @v1[dc] = 1.4
  print @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
  run
  alter @v1[dc] = 1.8
  print @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
  run
  alter @v1[dc] = 2
  print @m.xm1.msky130_fd_pr__nfet_01v8[vdsat]
  run

  plot (-dc1.i(v2)) (-dc2.i(v2)) (-dc3.i(v2)) (-dc4.i(v2)) (-dc5.i(v2))

.endc

.save all


 ** manual skywater pdks install (with patches applied)
* .lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /ef/tech/SW.2/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param mc_mm_switch=0
.param mc_pr_switch=0

**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
